module yArith(z,cout, a,b,ctrl);
 // add if ctrl =0, sub if ctrl =1
 output [31:0] z;
 output cout;
 input [31:0] a,b;
 input ctrl;
 wire [31:0] notB,tmp;
 wire cin;
 
 // instantiate compnents and connect them
 // just 4 lines of code
endmodule
